`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Hau Tao
//
// Create Date:    16:39:09 10/07/2015
// Module Name:    INCR
//////////////////////////////////////////////////////////////////////////////////
module INCR(pcout, pcin);

    input  [31:0] pcin;
    output [31:0] pcout;
    assign  pcout  = pcin + 1;

endmodule
