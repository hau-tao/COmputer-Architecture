
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Student: HAU TAO
// Create Date:    22:01:58 10/20/2015
// Module Name:    progrmCounter
//////////////////////////////////////////////////////////////////////////////////
module programCounter(npc, pc);
     input[31:0] npc;
     output [31:0] pc;
     assign pc = npc;
endmodule

